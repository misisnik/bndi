----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:22:41 11/12/2015 
-- Design Name: 
-- Module Name:    rom_1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity rom_4 is
    Port ( address : in  STD_LOGIC_VECTOR (12 downto 0);
           clk : in STD_LOGIC;
			  data: out  STD_LOGIC_VECTOR (3 downto 0));
end rom_4;

--rom 4 obsahuje 16bitove pismena a cisla
architecture Behavioral of rom_4 is
	--graphic database
	type rom_type is array(0 to 6655) of std_logic_vector(3 downto 0);
	constant database : rom_type :=
	(
		--cislo 0
		"1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0000", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "1011", 
		"1011", "1011", "0000", "0000", "0111", "0111", "0111", "0000", "0000", "0111", "0111", "0111", "0000", "0000", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "0000", "0000", "0111", "0111", "0111", "0000", "0000", "0111", "0111", "0111", "0000", "0000", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0000", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011",
		--cislo 1
		"1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0000", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011",
		--cislo 2
		"1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011",
		--cislo 3
		"1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011",
		--cislo 4
		"1011", "1011", "1011", "1011", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "1011", "1011",
		--cislo 5
		"1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011",
		--cislo 6
		"1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011",
		--cislo 7
		"1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011",
		--cislo 8
		"1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011",
		--cislo 9
		"1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011",
		---------
		--pismena a znaky
		---------
		--znak !
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011",
		--pismeno E
		"1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011",
		--pismeno T
		"1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011",
		--pismeno V
		"1011", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011",
		--pismeno Y
		"1011", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011",
		--pismeno P
		"1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011",
		--pismeno C
		"1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011",
		--pismeno D
		"1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011",
		--pismeno G
		"1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011",
		--pismeno A
		"1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0000", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "1011", 
		"1011", "1011", "0000", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0111", "0111", "0000", "0000", "1011", "1011", 
		"1011", "0000", "0000", "0111", "0111", "0000", "0000", "1011", "1011", "0000", "0000", "0111", "0111", "0000", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "1011", "1011", "1011", "1011", "0000", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "1011",
		--pismeno R
		"1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "1011", "1011",
		--pismeno M
		"1011", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0111", "0111", "0111", "0111", "0000", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "0000", "0111", "0111", "0000", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "0000", "0000", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "1011",
		--pismeno O
		"1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011",
		--pismeno X
		"1011", "1011", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0000", "1011", 
		"1011", "1011", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "1011", "1011",
		--pismeno S
		"1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "1011", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0111", "0111", "0111", "0000", "1011", 
		"1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", 
		"1011", "1011", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011",
		--button
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0000", "1011", "1011", "0000", "0000", "1011", "1011", "0000", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0000", "1011", "1011", "0000", "0000", "1011", "1011", "0000", "0000", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0000", "1011", "0000", "0000", "1011", "0000", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0100", "0100", "0100", "0100", "0100", "0100", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0100", "0100", "0100", "0100", "0100", "0100", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", 
		"1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", 
		"1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", 
		"1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011"
	);

begin
	process (clk)
	begin
		if (clk'event and clk = '1') then
			data <= database(to_integer(unsigned(address)));
		end if;
	end process;




end Behavioral;

