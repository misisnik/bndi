--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   15:26:31 10/26/2015
-- Design Name:   
-- Module Name:   C:/Users/xslade18/Desktop/bndi-master/keyboard_comunication/debouncer_test.vhd
-- Project Name:  keyboard_comunication
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: debouncer
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY debouncer_test IS
END debouncer_test;
 
ARCHITECTURE behavior OF debouncer_test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT debouncer
    PORT(
         clk : IN  std_logic;
         deb_in : IN  std_logic;
         deb_out : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal deb_in : std_logic := '0';

 	--Outputs
   signal deb_out : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: debouncer PORT MAP (
          clk => clk,
          deb_in => deb_in,
          deb_out => deb_out
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		
		deb_in <= '1';
		wait for 100 ns;
		deb_in <= '1';
		wait for 100 ns;
		deb_in <= '1';
		wait for 100 ns;
		deb_in <= '0';
		wait for 100 ns;
		deb_in <= '1';
		wait for 100 ns;
		deb_in <= '1';
		wait for 100 ns;
		
		deb_in <= '0';
		wait for 100 ns;
		deb_in <= '0';
		wait for 100 ns;
		deb_in <= '1';
		wait for 100 ns;
      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
