----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:22:41 11/12/2015 
-- Design Name: 
-- Module Name:    rom_1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity rom_1 is
    Port ( address : in  STD_LOGIC_VECTOR (14 downto 0);
           data : out  STD_LOGIC_VECTOR (3 downto 0));
end rom_1;

architecture Behavioral of rom_1 is
	--graphic database
	signal rom_data : std_logic_vector(3 downto 0);
	type rom_type is array(0 to 3071) of std_logic_vector(3 downto 0);
	constant database : rom_type :=
	(
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0010", "0010", "0010", "0010", "0010", "0000", "0000", "0000", "0000", "0000", "0010", "0010", "0010", "0010", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0010", "0010", "0010", "0010", "0000", "0111", "0111", "0111", "0111", "0111", "0000", "0010", "0010", "0010", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0010", "0010", "0010", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0010", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0010", "0010", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0010", "0010", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0010", "0010", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0010", "0010", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0010", "0010", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0010", "0010", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0010", "0010", "0010", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0110", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0010", "0010", "0010", "0000", "0111", "0111", "0111", "0111", "0111", "0000", "0110", "0110", "0110", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0010", "0000", "0000", "0000", "0000", "0000", "0110", "0110", "0110", "0110", "0110", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0100", "0100", "0100", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "0000", "0100", "0100", "0110", "0110", "0000", "0000", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0000", "0000", "0110", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "0000", "0100", "0100", "0000", "0110", "0110", "0110", "0000", "0000", "0110", "0110", "0110", "0110", "0110", "0000", "0000", "0110", "0110", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0100", "0100", "0000", "0000", "0000", "0110", "0110", "0110", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0110", "0110", "0110", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "0000", "0100", "0000", "0111", "0111", "0111", "0000", "0110", "0110", "0110", "0000", "0100", "0100", "0000", "0110", "0110", "0110", "0110", "0110", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0100", "0000", "0111", "0111", "0111", "0111", "0111", "0000", "0110", "0110", "0000", "0100", "0100", "0000", "0110", "0110", "0110", "0110", "0110", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "0000", "0100", "0000", "0111", "0111", "0111", "0111", "0111", "0000", "0110", "0110", "0110", "0000", "0000", "0110", "0110", "0110", "0110", "0110", "0110", "0000", "0111", "0111", "0111", "0000", "1011", "1011", "1011", "1011", 
		"1011", "1011", "0000", "0100", "0100", "0100", "0000", "0111", "0111", "0111", "0000", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0000", "0111", "0111", "0000", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "0000", "0100", "0100", "0100", "0100", "0000", "0000", "0000", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0000", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "0000", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0000", "0110", "0110", "0110", "0110", "0000", "0000", "0000", "0000", "0110", "0110", "0110", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"0000", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0000", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0000", "0110", "0110", "0110", "0110", "0110", "0110", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"0000", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0000", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0000", "0110", "0110", "0110", "0110", "0110", "0110", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011",
		--vrtula
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"0000", "0000", "1011", "1011", "1011", "1011", "0000", "0000", "1111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"0111", "0000", "0000", "1011", "1011", "0000", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"0111", "0000", "0000", "1011", "1011", "0000", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"0000", "0000", "1011", "1011", "1011", "1011", "0000", "0000", "1111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"0111", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"0000", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011",
		--vrtula2
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1111", "0000", "0000", "1011", "1011", "1011", "1011", "0000", "0000", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "0000", "0000", "0111", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0000", "0000", "1011", "1011", "0000", "0000", "0111", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1111", "0000", "0000", "1011", "1011", "1011", "1011", "0000", "0000", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1011", "1011", "1011", "1011", "1011", "1011", "0000", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", "0111", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0000", 
		"1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011"

	);
begin
	-- set data from database to output
	data <= database(to_integer(unsigned(address)));

end Behavioral;

